`timescale 1ns / 1ps

module DataMemory(input [31:0] mr, input [31:0] mqb, input mwmem, input clk, output reg [31:0] mdo);
    reg [31:0] memory [0:63];
    initial begin
        memory[0] = 'hA00000AA;
        memory[1] = 'h10000011;
        memory[2] = 'h20000022;
        memory[3] = 'h30000033;
        memory[4] = 'h40000044;
        memory[5] = 'h50000055;
        memory[6] = 'h60000066;
        memory[7] = 'h70000077;
        memory[8] = 'h80000088;
        memory[9] = 'h90000099;
    end
    always @ (*) begin
        mdo = memory[mr/4];
    end
    always @ (negedge clk) begin
        if(mwmem == 1) begin
            memory[mr] = mqb;
        end
    end
endmodule